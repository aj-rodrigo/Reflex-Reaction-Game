`timescale 1ns / 1ps

module Lights(rst, numIn, scoreIn, timerIn, sw, led);

input rst; 
input [4:0] numIn;
input [5:0] scoreIn, timerIn;
input [15:0] sw;
output [15:0] led;

reg [15:0] ledForm;


always @(*) begin
    if(rst)
        ledForm <= 16'b0000000000000010;
    else begin
        case(timerIn)
            30: ledForm <= 16'b1000000000000000;            //16'b1000000000000000;
            29: ledForm <= 16'b0010000000000000;            //16'b0100000000000000;
            28: ledForm <= 16'b0000000010000000;            //16'b0010000000000000;
            27: ledForm <= 16'b0000010000000000;            //16'b0001000000000000;
            26: ledForm <= 16'b0000001000000000;            //16'b0000100000000000;
            25: ledForm <= 16'b0000010000000000;            //16'b0000010000000000;
            24: ledForm <= 16'b0000001000000000;            //16'b0000001000000000;
            23: ledForm <= 16'b0000000100000000;            //16'b0000000100000000;
            22: ledForm <= 16'b0100000000000000;            //16'b0000000010000000;
            21: ledForm <= 16'b0000000000000100;            //16'b0000000001000000;
            20: ledForm <= 16'b0001000000000000;            //16'b0000000000100000;
            19: ledForm <= 16'b0000000000010000;            //16'b0000000000010000;
            18: ledForm <= 16'b0000001000000000;            //16'b0000000000001000;
            17: ledForm <= 16'b0000000000000100;            //16'b0000000000000100;
            16: ledForm <= 16'b0000000000000010;            //16'b0000000000000010;
            15: ledForm <= 16'b0000100000000000;            //16'b0000000000000001;
            14: ledForm <= 16'b0000000000000010;            //16'b0000000000000010;
            13: ledForm <= 16'b0000000100000000;            //16'b0000000000000100;
            12: ledForm <= 16'b0000000000001000;            //16'b0000000000001000;
            11: ledForm <= 16'b0000000000010000;            //16'b0000000000010000;
            10: ledForm <= 16'b0000000000100000;            //16'b0000000000100000;
            9:  ledForm <= 16'b0001000000000000;            //16'b0000000001000000;
            8:  ledForm <= 16'b0000000010000000;            //16'b0000000010000000;
            7:  ledForm <= 16'b0000000000010000;            //16'b0000000100000000;
            6:  ledForm <= 16'b0000001000000000;            //16'b0000001000000000;
            5:  ledForm <= 16'b0000010000000000;            //16'b0000010000000000;
            4:  ledForm <= 16'b0000100000000000;            //16'b0000100000000000;
            3:  ledForm <= 16'b0001000000000000;            //16'b0001000000000000;
            2:  ledForm <= 16'b0010000000000000;            //16'b0010000000000000;
            1:  ledForm <= 16'b0100000000000000;            //16'b0100000000000000;
            0:  ledForm <= 16'b1000000000000000;            //16'b1000000000000000;
        endcase
    end
end



assign led = ledForm;

endmodule
